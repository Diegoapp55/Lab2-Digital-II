`timescale 1ns / 1ps
module sh_r(
  input [2:0] portA,
  input init_sh_r,       //Pin para habilitar o no este módulo (Asignar a pulsador para que refresque y no se quede en 1)
  input clk,             //Pin para sincronizar con el reloj
  input rst,             //Pin para volver al dato sin corrimientos
  output [3:0] sal_sh_r  //Pines para extraer lo que retorna este módulo y usarlo en el top-module
);

reg [3:0] A; //Registro que almacenará el número desplazado
assign sal_sh_r = A;

always @ (posedge clk) begin
  if (rst) A = {1'b0,portA}; //Devuelve A a su posición original (En los últimos 3 LSB), es decir, reinicia el desplazamiento
  else if (init_sh_r) A <= A >> 1; //Desplaza A a la derecha
end

endmodule
